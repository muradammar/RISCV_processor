module datapath(

);

endmodule

